// set INCPHY_CELL    {FILLCAP3A10TR FILLCAP4A10TR FILLCAP8A10TR FILLCAP16A10TR FILLCAP32A10TR FILLCAP64A10TR FILLCAP128A10TR}
module FILLCAP3A10TR (); endmodule
module FILLCAP4A10TR (); endmodule
module FILLCAP8A10TR (); endmodule
module FILLCAP16A10TR (); endmodule
module FILLCAP32A10TR (); endmodule
module FILLCAP64A10TR (); endmodule
module FILLCAP128A10TR (); endmodule